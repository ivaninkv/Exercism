module main

fn color_code(color string) int {
	return colors.index(color)
}

const colors = ['black', 'brown', 'red', 'orange', 'yellow', 'green', 'blue', 'violet', 'grey',
	'white']
